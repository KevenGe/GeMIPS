/******************************************************************************
*   
*   文件名称：CTRL.v
*   文件说明：这个文件是GeMIPS的负责流水线暂停的模块。 
* 
*   作者：葛启丰
*   时间：2020-07-07
*
******************************************************************************/

module CTRL (

       );

endmodule
